module apb4_ps2 (
    input logic ps2_clk_i,
    input logic ps2_dat_i
);

endmodule

module ps2 ();
endmodule
