
module apb_timer (
    input logic clk,
    input logic rstn,
    input 
);
    
endmodule