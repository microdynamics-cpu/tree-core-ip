interface apb_if;
    
endinterface